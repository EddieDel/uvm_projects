`include "uvm_macros.svh"


package apb_test_pkg;
 import uvm_pkg::*;


 `include "apb_reg_model.sv";


endpackage
