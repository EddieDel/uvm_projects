`ifndef APB_ENV_PKG_SV
 `define APB_ENV_PKG_SV

`include "uvm_macros.svh"
`include "apb_agent_pkg.sv"
`include "apb_reg_pkg.sv"


package apb_env_pkg;
 import uvm_pkg::*;

 import apb_agent_pkg::*;
 import apb_reg_pkg::*;
 

 `include "apb_reg_adapter.sv";
 `include "apb_ral_sequences.sv";
 `include "apb_environment.sv";


endpackage
 

`endif
