`ifndef TEST_PKG_SV
 `define TEST_PKG_SV

`include "uvm_macros.svh"
`include "agent_pkg.sv"

package test_pkg;
import uvm_pkg::*;
import agent_pkg::*; 

`include "environment.sv";
 `include "test_base.sv";
 `include "test_counter.sv";
 


endpackage

`endif
